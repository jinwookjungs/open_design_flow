/home/jwjung/workspace/github/open_design_flow/bench/b19/b19.lef